module Instruction(clk,run,instruction,pc,addr_mem,addr_change);
input clk,run;
input [31:0]addr_change;

output [31:0] instruction;
output reg [29:0] pc=30'd0;

output wire [31:0] addr_mem;

reg [7:0] Mem [255:0];
integer i;
/*
initial
	for(i=0;i<256;i=i+1) Mem[i]<=i;*/
/*
initial
	begin
	Mem[0]  <=  32'b000000_00001_00010_00011_00000_100000;     //add   $3,$1,$2    3�żĴ���ֵΪ 3 
	Mem[1]  <=  32'b000000_00001_00010_00100_00000_100010;     //sub   $4,$1,$2    4�żĴ���ֵΪ -1
	Mem[2]  <=  32'b100011_00001_00101_00000_00000_000111;     //lw    $5,$1,7     5�żĴ���ֵΪ �洢�� 8
	Mem[3]  <=  32'b000000_00101_00001_00110_00000_100011;     //subu  $6,$5,$1    6�żĴ���ֵΪ 8-1=7
	Mem[4]  <=  32'b000100_00001_00001_00000_00000_000010;     //beq   $1,$1,2      PC+1+2=4+1+2=7, ��һ����PC=7     4
	Mem[5]  <=  32'b000000_00001_00010_00101_00000_101011;
	Mem[6]  <=  32'b101011_00001_00011_00000_00000_000101;
	Mem[7]  <=  32'b000000_00100_00001_00111_00000_101010;      //slt   $7,$4,$1    �з���С����1    7�żĴ���ֵΪ 1
	Mem[8]  <=  32'b000000_00100_00001_01000_00000_101011;      //sltu  $8,$4,$1    �޷���С����1    8�żĴ���ֵΪ 0
	Mem[9]  <=  32'b001001_00001_01001_11111_11111_111000;      //addiu $9, $1,������
	Mem[10]  <=  32'b101011_00001_01010_00000_00000_001111;      //sw    $10,$1,15   ��10�żĴ�����ֵ�浽 �洢�� 16��
	Mem[11]  <=  32'b001101_00111_01011_00000_00000_000010;      //ori   $11,$7,2   7�żĴ���ֵΪ 1 ��2  ���,���Ϊ3 ��11�żĴ���
	Mem[12]  <=  32'b000010_00000_00000_00000_00000_000010;      //jump  ��תָ�   ��ת��14
	end*/

initial
	begin
	{Mem[0],Mem[1],Mem[2],Mem[3]}      <=  32'b000000_00001_00010_00011_00000_100000;     //add   $3,$1,$2    3�żĴ���ֵΪ 3 
	{Mem[4],Mem[5],Mem[6],Mem[7]}      <=  32'b000000_00001_00010_00100_00000_100010;     //sub   $4,$1,$2    4�żĴ���ֵΪ -1
	{Mem[8],Mem[9],Mem[10],Mem[11]}    <=  32'b100011_00001_00101_00000_00000_000111;     //lw    $5,$1,7     5�żĴ���ֵΪ �洢�� 8
	{Mem[12],Mem[13],Mem[14],Mem[15]}  <=  32'b000000_00101_00001_00110_00000_100011;     //subu  $6,$5,$1    6�żĴ���ֵΪ 8-1=7
	{Mem[16],Mem[17],Mem[18],Mem[19]}  <=  32'b000100_00001_00001_00000_00000_000010;     //beq   $1,$1,2      PC+1+2=4+1+2=7, ��һ����PC=7     4
	{Mem[20],Mem[21],Mem[22],Mem[23]}  <=  32'b000000_00001_00010_00101_00000_101011;	//sltu $5,$1,$2  �޷���С����1    5�żĴ���ֵΪ 1
	{Mem[24],Mem[25],Mem[26],Mem[27]}  <=  32'b101011_00001_00011_00000_00000_000101;	//sw $3,$1,5    ��3�żĴ�����ֵ�浽 �洢�� 6��
	{Mem[28],Mem[29],Mem[30],Mem[31]}  <=  32'b000000_00100_00001_00111_00000_101010;      //slt   $7,$4,$1    �з���С����1    7�żĴ���ֵΪ 1
	{Mem[32],Mem[33],Mem[34],Mem[35]}  <=  32'b000000_00100_00001_01000_00000_101011;      //sltu  $8,$4,$1    �޷���С����1    8�żĴ���ֵΪ 0
	{Mem[36],Mem[37],Mem[38],Mem[39]}  <=  32'b001001_00001_01001_11111_11111_111000;      //addiu $9, $1,������
	{Mem[40],Mem[41],Mem[42],Mem[43]}  <=  32'b101011_00001_01010_00000_00000_001111;      //sw    $10,$1,15   ��10�żĴ�����ֵ�浽 �洢�� 16��
	{Mem[44],Mem[45],Mem[46],Mem[47]}  <=  32'b001101_00111_01011_00000_00000_000010;      //ori   $11,$7,2   7�żĴ���ֵΪ 1 ��2  ���,���Ϊ3 ��11�żĴ���
	{Mem[48],Mem[49],Mem[50],Mem[51]}  <=  32'b000010_00000_00000_00000_00000_000010;      //jump  ��תָ�   ��ת��2
	end
/*
always@(*)
begin
	Mem[0] =8'b0000_0000; Mem[1] =8'b0010_0010;  Mem[2] =8'b0001_1000; Mem[3] =8'b0010_0000;//add   $3,$1,$2    3�żĴ���ֵΪ 3
	Mem[4] =8'b0000_0000; Mem[5] =8'b0010_0010;  Mem[6] =8'b0010_0000; Mem[7] =8'b0010_0010;//sub   $4,$1,$2    4�żĴ���ֵΪ -1
	Mem[8] =8'b1000_1100; Mem[9] =8'b0010_0101;  Mem[10]=8'b0000_0000; Mem[11]=8'b0000_0111; //lw  $5,$1,7
	Mem[12]=8'b0000_0000; Mem[13]=8'b1010_0001;  Mem[14]=8'b0011_0000; Mem[15]=8'b0010_0011;//subu  $6,$5,$1    6�żĴ���ֵΪ 8-1=7
	Mem[16]=8'b0001_0000; Mem[17]=8'b0010_0001;  Mem[18]=8'b0000_0000; Mem[19]=8'b0000_0010;//beq   $1,$1,2      PC+1+2=4+1+2=7, ��һ����PC=7     4
	Mem[20]=8'b0000_0000; Mem[21]=8'b0010_0010;  Mem[22]=8'b0010_1000; Mem[23]=8'b0010_1011;//sltu $5,$1,$2  �޷���С����1    5�żĴ���ֵΪ 1
	Mem[24]=8'b1010_1100; Mem[25]=8'b0010_0011;  Mem[26]=8'b0000_0000; Mem[27]=8'b0000_0101;//sw $3,$1,5    ��3�żĴ�����ֵ�浽 �洢�� 6��
	Mem[28]=8'b0000_0000; Mem[29]=8'b1000_0001;  Mem[30]=8'b0011_1000; Mem[31]=8'b0010_1010;//slt   $7,$4,$1    �з���С����1    7�żĴ���ֵΪ 1
	Mem[32]=8'b0000_0000; Mem[33]=8'b1000_0001;  Mem[34]=8'b0100_0000; Mem[35]=8'b0010_1011;//sltu  $8,$4,$1    �޷���С����1    8�żĴ���ֵΪ 0
	Mem[36]=8'b0010_0100; Mem[37]=8'b0010_1001;  Mem[38]=8'b1111_1111; Mem[39]=8'b1111_1000;//addiu $9, $1,������
	Mem[40]=8'b1010_1100; Mem[41]=8'b0010_1010;  Mem[42]=8'b0000_0000; Mem[43]=8'b0000_1111;//sw    $10,$1,15   ��10�żĴ�����ֵ�浽 �洢�� 16��
	Mem[44]=8'b0011_0100; Mem[45]=8'b1110_1011;  Mem[46]=8'b0000_0000; Mem[47]=8'b0000_0010;//ori   $11,$7,2   7�żĴ���ֵΪ 1 ��2  ���,���Ϊ3 ��11�żĴ���
	Mem[48] =8'b0000_0000; Mem[49] =8'b0010_1011;  Mem[50] =8'b0010_1000; Mem[51] =8'b0010_0000; //add $5,$1,$11
	Mem[52]=8'b0000_1000; Mem[53]=8'b0000_0000;  Mem[54]=8'b0000_0000; Mem[55]=8'b0000_0010;//jump  ��תָ�   ��ת��2
	instruction={Mem[addr_mem],Mem[addr_mem+1],Mem[addr_mem+2],Mem[addr_mem+3]};
end*/

//assign instruction={Mem[addr_mem],Mem[addr_mem+1],Mem[addr_mem+2],Mem[addr_mem+3]};

wire [29:0]temp1;
wire [29:0]temp2;
reg [29:0]temp3;
reg [31:0]temp4;
wire [29:0]M2;
assign instruction={Mem[addr_mem],Mem[addr_mem+1],Mem[addr_mem+2],Mem[addr_mem+3]};
assign temp1=pc;
assign temp2=instruction[15:0];
assign addr_mem = (addr_change==32'b0)?temp4:addr_change;
always@(negedge clk)
begin 
	/*
	pc=temp4[31:2];
	temp3 = pc + 1 + (branch_zero ? instruction[15:0] : 0);
	temp4 ={(jump?M2:temp3),2'b00};
	*/
	
	//ֻ��PC+1,run=0ʱpc����
	if(run==0)
	begin
		pc=addr_mem[31:2];
		pc=pc+1;
		temp4={pc,2'b00};
	end
end
//mux2to1 mux1(clk,temp1,temp2,branch_zero,temp3); // branch  ��ת��ַ
//assign temp3 = temp1 + 1 + (branch_zero ? temp2 : 0);


//assign M2={pc[29:26],instruction[25:0]};          // jump    ��ת��ַ


//mux2to1_29 mux2(clk,temp3,M2,jump,temp4);
//assign temp4={(jump?M2:temp3),2'b00};

endmodule